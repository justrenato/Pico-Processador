entity test is
end test;
